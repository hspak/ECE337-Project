// $Id: $
// File name:   fader_wrapper.sv
// Created:     4/23/2014
// Author:      Patrick Gohier
// Lab Section: 337-04
// Version:     1.0  Initial Design Entry
// Description: Fader Multiplier Wrapper
module fader_wrapper (
  
);

endmodule
